class pkt1;
    string mode;

endclass //pkt1